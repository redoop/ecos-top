`timescale 1ns / 1ps

module soc_tb ();
  localparam real OSC_CLK_25M_PEROID = 40;

  wire ext_rst_n_i_pad;
  wire osc_clk_25m_i_pad;
  wire old_ip_spi_flash_clk_pad;
  wire [1:0] old_ip_spi_flash_cs_pad;
  wire old_ip_spi_flash_mosi_pad;
  wire old_ip_spi_flash_miso_pad;
  wire old_ip_uart_rx_pad;
  wire old_ip_uart_tx_pad;

  logic r_osc_clk_25m, r_ext_rst_n;
  logic [2:0] r_ip_sel;

  assign osc_clk_25m_i_pad = r_osc_clk_25m;
  assign ext_rst_n_i_pad = r_ext_rst_n;

  asic_top u_asic_top (
      .ip_sel_pad0       (r_ip_sel[0]),
      .ip_sel_pad1       (r_ip_sel[1]),
      .ip_sel_pad2       (r_ip_sel[2]),
      .sys_clk_i_pad     (osc_clk_25m_i_pad),
      .sys_clk_o_pad     (),
      .rst_n_pad         (ext_rst_n_i_pad),
      .io_pad0           (old_ip_uart_rx_pad),
      .io_pad1           (old_ip_uart_tx_pad),
      .io_pad2           (old_ip_spi_flash_clk_pad),
      .io_pad3           (old_ip_spi_flash_cs_pad[0]),
      .io_pad4           (old_ip_spi_flash_cs_pad[1]),
      .io_pad5           (),
      .io_pad6           (),
      .io_pad7           (),
      .io_pad8           (),
      .io_pad9           (),
      .io_pad10          (),
      .io_pad11          (old_ip_spi_flash_mosi_pad),
      .io_pad12          (old_ip_spi_flash_miso_pad),
      .io_pad13          (1'b0),
      .io_pad14          (1'b0),
      .io_pad15          (1'b0),
      .io_pad16          (),
      .io_pad17          (),
      .io_pad18          (),
      .io_pad19          (),
      .io_pad20          (),
      .io_pad21          (),
      .io_pad22          (),
      .io_pad23          (),
      .io_pad24          (),
      .io_pad25          (),
      .io_pad26          (),
      .io_pad27          (),
      .io_pad28          (),
      .io_pad29          (),
      .io_pad30          (),
      .io_pad31          (),
      .io_pad32          (),
      .io_pad33          (),
      .io_pad34          (),
      .io_pad35          (),
      .io_pad36          (),
      .io_pad37          (),
      .io_pad38          (),
      .io_pad39          (),
      .io_pad40          (),
      .io_pad41          (),
      .io_pad42          (),
      .io_pad43          (),
      .io_pad44          (),
      .io_pad45          (),
      .io_pad46          (),
      .io_pad47          (),
      .io_pad48          (),
      .io_pad49          (),
      .io_pad50          (),
      .io_pad51          (),
      .io_pad52          (),
      .io_pad53          (),
      .io_pad54          (),
      .io_pad55          (),
      .io_pad56          (),
      .io_pad57          (),
      .io_pad58          (),
      .io_pad59          (),
      .io_pad60          (),
      .io_pad61          (),
      .io_pad62          (),
      .io_pad63          (),
      .io_pad64          (),
      .io_pad65          (),
      .io_pad66          (),
      .io_pad67          (),
      .io_pad68          (),
      .io_pad69          (),
      .io_pad70          (),
      .io_pad71          (),
      .io_pad72          (),
      .io_pad73          (),
      .io_pad74          (),
      .io_pad75          (),
      .io_pad76          (),
      .io_pad77          (),
      .io_pad78          (),
      .io_pad79          (),
      .io_pad80          (),
      .io_pad81          ()
  );

  N25Qxxx u_old_ip_spi_N25Qxxx (
      .C_       (old_ip_spi_flash_clk_pad),
      .S        (old_ip_spi_flash_cs_pad[0]),
      .DQ0      (old_ip_spi_flash_mosi_pad),
      .DQ1      (old_ip_spi_flash_miso_pad),
      .HOLD_DQ3 (),
      .Vpp_W_DQ2(),
      .Vcc      ('d3000)
  );

  tty #(115200, 0) u_old_ip_uart_tty (
      .STX(old_ip_uart_rx_pad),
      .SRX(old_ip_uart_tx_pad)
  );

  task sim_reset(int delay);
    r_ext_rst_n = 1'b0;
    repeat (delay) @(posedge osc_clk_25m_i_pad);
    #1 r_ext_rst_n = 1'b1;
  endtask

  initial begin
    r_osc_clk_25m = 1'b0;
    forever begin
      #(OSC_CLK_25M_PEROID / 2) r_osc_clk_25m <= ~r_osc_clk_25m;
    end
  end
    
  // BitNet加速器测试激励
  initial begin
    // 等待复位完成
    wait(r_ext_rst_n == 1'b1);
    repeat(100) @(posedge osc_clk_25m_i_pad);
    
    $display("[%0t] Starting BitNet & Compact Accelerator Interface Test", $time);
    
    // 选择IP1 (SimpleEdgeAiSoC) - BitNet加速器
    r_ip_sel = 3'd1;
    repeat(100) @(posedge osc_clk_25m_i_pad);
    
    $display("[%0t] IP1 selected, BitNet & Compact SoC active with new interfaces", $time);
    
    // 等待系统完全稳定
    repeat(10000) @(posedge osc_clk_25m_i_pad);
    
    // 这里可以添加更多具体的BitNet和Compact接口测试
    $display("[%0t] BitNet & Compact interface signals now connected to asic_top", $time);
    
    // 运行一段时间让加速器处理数据
    repeat(100000) @(posedge osc_clk_25m_i_pad);
    
    $display("[%0t] BitNet & Compact Accelerator Interface Test Phase Completed", $time);
  end

  // BitNet加速器测试任务
  task test_bitnet_accel();
    // 等待复位完成
    wait(r_ext_rst_n == 1'b1);
    repeat(100) @(posedge osc_clk_25m_i_pad);
    
    $display("[%0t] Starting BitNet Accelerator Test", $time);
    
    // 选择IP1 (SimpleEdgeAiSoC)
    r_ip_sel = 3'd1;
    repeat(10) @(posedge osc_clk_25m_i_pad);
    
    // 等待系统稳定
    repeat(1000) @(posedge osc_clk_25m_i_pad);
    
    $display("[%0t] BitNet Accelerator Test Completed", $time);
  endtask

  // RISC-V 功能测试任务
  task test_riscv_functionality();
    reg [31:0] prev_gpio, curr_gpio;
    reg activity_detected;
    integer test_cycles;
    
    $display("[%0t] Starting RISC-V Core Functionality Test", $time);
    
    // 监控 GPIO 输出变化 (表明 CPU 活动)
    prev_gpio = u_asic_top.ip1_io_gpio_out;
    activity_detected = 1'b0;
    test_cycles = 0;
    
    repeat(10000) begin
      @(posedge osc_clk_25m_i_pad);
      curr_gpio = u_asic_top.ip1_io_gpio_out;
      test_cycles = test_cycles + 1;
      
      if (curr_gpio !== prev_gpio) begin
        activity_detected = 1'b1;
        $display("[%0t] RISC-V activity detected - GPIO changed: 0x%08x -> 0x%08x", 
                 $time, prev_gpio, curr_gpio);
        break;
      end
      
      // 检查异常信号
      if (u_asic_top.ip1_io_trap == 1'b1) begin
        $display("[%0t] RISC-V trap signal detected", $time);
      end
      
      // 检查中断信号
      if (u_asic_top.ip1_io_uart_tx_irq || u_asic_top.ip1_io_uart_rx_irq) begin
        $display("[%0t] UART interrupt detected", $time);
      end
    end
    
    if (activity_detected) begin
      $display("[%0t] ✅ RISC-V Core Test PASSED - CPU activity confirmed", $time);
    end else begin
      $display("[%0t] ⚠️  RISC-V Core Test - No GPIO activity (may be normal)", $time);
    end
    
    $display("[%0t] RISC-V test cycles completed: %0d", $time, test_cycles);
  endtask

  initial begin
      sim_reset(400);
      
      // 启动RISC-V功能测试
      test_riscv_functionality();
      
      // 启动BitNet测试
      test_bitnet_accel();
      
      // 运行足够长时间观察结果
      #50000000;
      
      $display("[%0t] All tests completed", $time);
      $finish;
  end

    initial begin
        if      ($test$plusargs("ip_sel00")) r_ip_sel = 3'd0;
        else if ($test$plusargs("ip_sel01")) r_ip_sel = 3'd1;
        else if ($test$plusargs("ip_sel02")) r_ip_sel = 3'd2;
        else if ($test$plusargs("ip_sel03")) r_ip_sel = 3'd3;
        else if ($test$plusargs("ip_sel04")) r_ip_sel = 3'd4;
        else if ($test$plusargs("ip_sel05")) r_ip_sel = 3'd5;

        if ($test$plusargs("dump_all")) begin
          $fsdbDumpfile("soc_tb.fsdb");
          $fsdbDumpvars(0, soc_tb, "+all");
        end

`ifdef VCD_DUMP
        // VCD dump for GTKWave
        $dumpfile("soc_tb.vcd");
        $dumpvars(0, soc_tb);
`endif

        if      ($test$plusargs("asm-flash"))       #1000000    $finish;
        else if ($test$plusargs("hello-flash"))     #1000000    $finish;
        else if ($test$plusargs("hello-mem"))     #40000000   $finish;
        else if ($test$plusargs("hello-sdram"))   #40000000   $finish;
        else if ($test$plusargs("memtest-flash"))   #600000000  $finish;
        else if ($test$plusargs("memtest-mem"))     #120000000  $finish;
        else if ($test$plusargs("memtest-sdram")) #60000000   $finish;
        else if ($test$plusargs("rtthread-flash"))  #1600000000 $finish;
        else if ($test$plusargs("rtthread-mem"))    #200000000  $finish;
        else if ($test$plusargs("rtthread-sdram"))  #200000000  $finish;
        else if ($test$plusargs("bitnet-test"))     #100000000  $finish;

    end

endmodule